module AXI_Interface (
    
);

//AXI����ģ�� ������AXI�ӿڷ������������/�����źŵ�

endmodule //AXI_Interface