module DCache(
    
);

endmodule //DCache