`ifndef AXICACHE_DEFINES_VH
    `define AXICACHE_DEFINES_VH

`endif 