`include "global_defines.vh"

module ITLB_stage(
    input         clk,
    input         reset,
    input             ITLB_found,
    input      [31:0] ITLB_VAddr, //���ַ
    output reg [31:0] ITLB_RAddr, //ʵ��ַ
    input      [ 3:0] ITLB_index,
    input      [19:0] ITLB_pfn,
    input      [ 3:0] ITLB_asid, //ASID
    input      [ 2:0] ITLB_c,
    input             ITLB_d,
    input             ITLB_v,
    output reg        ITLB_EX_Refill,
    output reg        ITLB_EX_Invalid //
);

always @(*) begin
    if(ITLB_VAddr[31:28] == 4'hA || ITLB_VAddr[31:28] == 4'hB) //ʵ��ַ�������λ����
        ITLB_RAddr <= {3'b000, ITLB_VAddr[28:0]};
    else if(ITLB_VAddr[31:28] == 4'h8 || ITLB_VAddr[31:28] == 4'h9) //ʵ��ַ�����λ����
        ITLB_RAddr <= {1'b0  , ITLB_VAddr[30:0]};
    else
        ITLB_RAddr <= {ITLB_pfn,ITLB_VAddr[11:0]};
end

always @(*) begin
    if(~ITLB_found && (ITLB_VAddr[31:28] <= 4'h7 || ITLB_VAddr[31:28] >= 4'hC))
        ITLB_EX_Refill <= 1'b1;
    else
        ITLB_EX_Refill <= 1'b0;
end

always @(*) begin
    if(ITLB_found && (ITLB_VAddr[31:28] <= 4'h7 || ITLB_VAddr[31:28] >= 4'hC) && ~ITLB_v)
        ITLB_EX_Invalid <= 1'b1;
    else
        ITLB_EX_Invalid <= 1'b0;
end

reg ITLB_Buffer_Hit;
wire ITLB_Buffer_valid;
always @(*) begin
    if(ITLB_VAddr[31:28] < 4'hC && ITLB_VAddr[31:28] > 4'h7)
        ITLB_Buffer_Hit = 1'b1;
    else if(ITLB_VAddr[31:13] == ITLB_pfn && ITLB_Buffer_valid)
        ITLB_Buffer_Hit = 1'b1;
    else 
        ITLB_Buffer_Hit = 1'b0;
end


parameter   IDLE =   4'd0,
            SEARCH = 4'd1;
reg ITLB_cstate;
reg ITLB_nstate;  
wire ITLB_Buffer_Wr;

always @(posedge clk) begin
    if(reset) begin
        ITLB_cstate <= IDLE;
    end else begin
        ITLB_cstate <= ITLB_nstate;
    end    
end

always @(*) begin
        case(ITLB_cstate)
            IDLE :
               if(ITLB_Buffer_Hit == 1'b0) begin
                    ITLB_nstate = SEARCH;
                end
                else begin
                   ITLB_nstate = IDLE;
                end
            SEARCH :
                 if(ITLB_Buffer_Hit == 1'b1) begin
                    ITLB_nstate = IDLE;
                end  
                else begin
                    ITLB_nstate = SEARCH; 
                end         
     endcase
end

assign ITLB_Buffer_Wr  = (ITLB_cstate == SEARCH);  //��state2״̬�´�TLB Buffer��дʹ��
endmodule