module regfile(
    input         clk,
    input         reset,
    // READ PORT 1
    input  [ 4:0] raddr1,
    output [31:0] rdata1,
    // READ PORT 2
    input  [ 4:0] raddr2,
    output [31:0] rdata2,
    // WRITE PORT
    input         we,       //write enable, HIGH valid
    input  [ 4:0] waddr,
    input  [31:0] wdata,
    output [31:0] stack_addr
);
reg [31:0] rf[31:0];

assign stack_addr = rf[31];

integer i;
//WRITE
always @(posedge clk) begin
    if(reset) begin
        for (i = 0; i < 6'd32; i = i + 1) begin
            rf[i] <= 32'b0;
        end
    end
    else if (we) rf[waddr]<= wdata;
end

//READ OUT 1
assign rdata1 = (raddr1==5'b0) ? 32'b0 : rf[raddr1];

//READ OUT 2
assign rdata2 = (raddr2==5'b0) ? 32'b0 : rf[raddr2];

endmodule