`include "global_defines.vh"

module BPU#(
    parameter  DATA_WIDTH       =   64, // 前两位是饱和计数器，中间22位是tag，后32位是目标地址
    parameter  PHT_NUMS         =   256,
    parameter  W_Taken          =   2'b00,
    parameter  S_Taken          =   2'b01,
    parameter  WN_Taken         =   2'b10,
    parameter  SN_Taken         =   2'b11
)
(
    input clk,
    input reset,
    input [31:0] fs_pc,//连temp_fs_pc
    input ds_allowin,
    input [`BRESULT_WD - 1 :0] BResult,
    output [31:0] target,
    output BPU_valid,
    output [`BPU_TO_DS_BUS_WD-1:0] BPU_to_ds_bus
);
reg [7:0] BHR_cnt;
/*************************写入PHT*************************************/
reg [31:0] BPU_es_pc;
reg [1:0] BPU_old_Count;
reg BPU_is_branch;
//reg BPU_br_stall;
reg BPU_br_taken;
reg [31:0] BPU_br_target;
reg [3:0] branch_type;
always @(posedge clk) begin
    {   branch_type,
        BHR_cnt,
        BPU_es_pc,      //跳转指令的PC
        BPU_old_Count,  //跳转指令PC跳转次数的历史记录，2位饱和计数器，需更新后再写入PHT
        BPU_is_branch,  //PC是否是跳转指令
        //BPU_br_stall,  // 当判断阶段已到exe阶段时，此信号可删除
        BPU_br_taken,   //是否成功跳转
        BPU_br_target   //跳转的目标地址
                        } <=  BResult;
end

wire PHT_we;
wire [7:0] PHT_wr_index;
wire [21:0] PHT_wr_tag;
reg [1:0] BPU_new_Count;
wire [DATA_WIDTH-1 : 0] PHT_wr_data;//根据BResult得出

always @(*) begin
    if(BHR_cnt[2:0]==BHR_cnt[5:3]&& ((branch_type==`BRANCH_TYPE_BEQ) 
    || (branch_type==`BRANCH_TYPE_BNE)  || (branch_type==`BRANCH_TYPE_BGEZ) 
    || (branch_type==`BRANCH_TYPE_BGTZ) || (branch_type==`BRANCH_TYPE_BLEZ) 
    || (branch_type==`BRANCH_TYPE_BLTZ) || (branch_type==`BRANCH_TYPE_BGEZAL) 
    || (branch_type==`BRANCH_TYPE_BLTZAL) ))
        BPU_new_Count = {2{BHR_cnt[2]}} ;
    else if(BHR_cnt[3:0]==BHR_cnt[7:4]&& ((branch_type==`BRANCH_TYPE_BEQ) 
    || (branch_type==`BRANCH_TYPE_BNE)  || (branch_type==`BRANCH_TYPE_BGEZ) 
    || (branch_type==`BRANCH_TYPE_BGTZ) || (branch_type==`BRANCH_TYPE_BLEZ) 
    || (branch_type==`BRANCH_TYPE_BLTZ) || (branch_type==`BRANCH_TYPE_BGEZAL) 
    || (branch_type==`BRANCH_TYPE_BLTZAL) ))
        BPU_new_Count = {2{BHR_cnt[3]}} ;
    else if(BHR_cnt[2:0]==BHR_cnt[7:5]&& ((branch_type==`BRANCH_TYPE_BEQ) 
    || (branch_type==`BRANCH_TYPE_BNE)  || (branch_type==`BRANCH_TYPE_BGEZ) 
    || (branch_type==`BRANCH_TYPE_BGTZ) || (branch_type==`BRANCH_TYPE_BLEZ) 
    || (branch_type==`BRANCH_TYPE_BLTZ) || (branch_type==`BRANCH_TYPE_BGEZAL) 
    || (branch_type==`BRANCH_TYPE_BLTZAL) ))
        BPU_new_Count = {2{BHR_cnt[3]}} ; 
    else if(BHR_cnt[1:0]==BHR_cnt[7:6]&& ((branch_type==`BRANCH_TYPE_BEQ) 
    || (branch_type==`BRANCH_TYPE_BNE)  || (branch_type==`BRANCH_TYPE_BGEZ) 
    || (branch_type==`BRANCH_TYPE_BGTZ) || (branch_type==`BRANCH_TYPE_BLEZ) 
    || (branch_type==`BRANCH_TYPE_BLTZ) || (branch_type==`BRANCH_TYPE_BGEZAL) 
    || (branch_type==`BRANCH_TYPE_BLTZAL) ))
        BPU_new_Count = {2{BHR_cnt[2]}} ;    
    // if(BHR_cnt[3:0]==4'b1111 && ((branch_type==`BRANCH_TYPE_BEQ) 
    // || (branch_type==`BRANCH_TYPE_BNE)  || (branch_type==`BRANCH_TYPE_BGEZ) 
    // || (branch_type==`BRANCH_TYPE_BGTZ) || (branch_type==`BRANCH_TYPE_BLEZ) 
    // || (branch_type==`BRANCH_TYPE_BLTZ) || (branch_type==`BRANCH_TYPE_BGEZAL) 
    // || (branch_type==`BRANCH_TYPE_BLTZAL) ))
    //     BPU_new_Count = S_Taken ;
    // else if(BHR_cnt[3:0]==4'b0111  && ((branch_type==`BRANCH_TYPE_BEQ) 
    // || (branch_type==`BRANCH_TYPE_BNE)  || (branch_type==`BRANCH_TYPE_BGEZ) 
    // || (branch_type==`BRANCH_TYPE_BGTZ) || (branch_type==`BRANCH_TYPE_BLEZ) 
    // || (branch_type==`BRANCH_TYPE_BLTZ) || (branch_type==`BRANCH_TYPE_BGEZAL) 
    // || (branch_type==`BRANCH_TYPE_BLTZAL) ) )
    //     BPU_new_Count = {2{BHR_cnt[4]}} ;
    // else if(BHR_cnt[3:0]==4'b1000  && ((branch_type==`BRANCH_TYPE_BEQ) 
    // || (branch_type==`BRANCH_TYPE_BNE)  || (branch_type==`BRANCH_TYPE_BGEZ) 
    // || (branch_type==`BRANCH_TYPE_BGTZ) || (branch_type==`BRANCH_TYPE_BLEZ) 
    // || (branch_type==`BRANCH_TYPE_BLTZ) || (branch_type==`BRANCH_TYPE_BGEZAL) 
    // || (branch_type==`BRANCH_TYPE_BLTZAL) ))
    //     BPU_new_Count = {2{BHR_cnt[4]}} ;
    // else if(BHR_cnt[3:0]==4'b0000   && ((branch_type==`BRANCH_TYPE_BEQ) 
    // || (branch_type==`BRANCH_TYPE_BNE)  || (branch_type==`BRANCH_TYPE_BGEZ) 
    // || (branch_type==`BRANCH_TYPE_BGTZ) || (branch_type==`BRANCH_TYPE_BLEZ) 
    // || (branch_type==`BRANCH_TYPE_BLTZ) || (branch_type==`BRANCH_TYPE_BGEZAL) 
    // || (branch_type==`BRANCH_TYPE_BLTZAL) ))
    //     BPU_new_Count = SN_Taken ;
    // else 
        case (BPU_old_Count)
            SN_Taken: BPU_new_Count = BPU_br_taken ? WN_Taken : SN_Taken;
            WN_Taken: BPU_new_Count = BPU_br_taken ? W_Taken  : SN_Taken;
            W_Taken : BPU_new_Count = BPU_br_taken ? S_Taken  : WN_Taken;
            S_Taken : BPU_new_Count = BPU_br_taken ? W_Taken  : S_Taken;    
            default: BPU_new_Count = W_Taken;
        endcase
end

assign PHT_we = BPU_is_branch;
assign PHT_wr_index = BPU_es_pc[9:2] ;
assign PHT_wr_tag = BPU_es_pc[31:10];
assign PHT_wr_data = {BHR_cnt,BPU_new_Count, PHT_wr_tag, BPU_br_target};

/*************************************************************************/

/*****************************读PHT***********************************/

wire [7:0] PHT_rd_index;      //读地址
wire [21:0] PHT_rout_tag;      //读出的tag
wire [31:0] PHT_rout_target;   //读出的目标地址
wire [1:0] PHT_rout_Count;    //读出的饱和计数器
wire [7:0] BHR_rout_cnt;
wire PHT_hit;
wire [DATA_WIDTH-1 : 0] PHT_rd_data;//读出的PHT
assign PHT_rd_index = fs_pc[9:2] ;
assign {BHR_rout_cnt,PHT_rout_Count,PHT_rout_tag,PHT_rout_target} = PHT_rd_data;
assign PHT_hit  = (PHT_rout_tag == fs_pc[31:10]) & ~PHT_we; // 写的时候返回数据不是想要读的

wire [21:0] debug_fs_pc_tag;
assign debug_fs_pc_tag = fs_pc[31:10];


wire [31:0] BPU_ret_addr;

reg BPU_valid_reg;
reg [31:0] BPU_ret_addr_reg;
reg [1:0] BPU_Count_reg;
reg BPU_is_taken_reg;               //预测是否跳转
reg [7:0] BHR_cnt_reg;
//reg [3:0]branch_type;
assign BPU_to_ds_bus = {
                            BHR_cnt_reg,   
                            BPU_is_taken_reg,
                            BPU_Count_reg,
                            BPU_valid_reg,
                            BPU_ret_addr_reg
                            };
assign BPU_ret_addr = PHT_rout_Count[1] ? fs_pc + 8 : PHT_rout_target;
// always @(posedge clk) begin
//     if(reset)begin
//         branch_type <=0;
//     end
//     else begin
//         branch_type <= branch_type;
//     end
//end 

always @(posedge clk) begin
    if(reset)begin
        BPU_valid_reg <= 0;
        BPU_Count_reg <= 0;
        BPU_ret_addr_reg <= 0;
        BPU_is_taken_reg <= 0;
        BHR_cnt_reg  <=0;
    end

    if(ds_allowin)begin
        if(PHT_hit)begin
            BPU_valid_reg <= 1;
            BPU_Count_reg <= PHT_rout_Count;
            BPU_ret_addr_reg <= BPU_ret_addr;
            BPU_is_taken_reg <= ~PHT_rout_Count[1];
            BHR_cnt_reg <= BHR_rout_cnt;
        end
        else begin
            BPU_valid_reg <= 0;
           // BPU_Count_reg <= 0;
            BPU_ret_addr_reg <= 0;
            BPU_is_taken_reg <= 0;
            BHR_cnt_reg  <=0;
        end
    end
    
end

/*************************************************************************/

/*****************************BHR*****************************************/

always @(posedge clk) begin
    if(reset) begin
        BHR_cnt <= 0;
    end
    else if(PHT_we &&  ((branch_type==`BRANCH_TYPE_BEQ) 
    || (branch_type==`BRANCH_TYPE_BNE)  || (branch_type==`BRANCH_TYPE_BGEZ) 
    || (branch_type==`BRANCH_TYPE_BGTZ) || (branch_type==`BRANCH_TYPE_BLEZ) 
    || (branch_type==`BRANCH_TYPE_BLTZ) || (branch_type==`BRANCH_TYPE_BGEZAL) 
    || (branch_type==`BRANCH_TYPE_BLTZAL) )) begin
        BHR_cnt <= {BHR_cnt[6:0],BPU_br_taken};
        end
    else begin
        BHR_cnt <= BHR_cnt;
    end
    
end
    
/*************************************************************************/

assign target = BPU_ret_addr;
assign BPU_valid = PHT_hit;
assign Count = BPU_Count_reg;

wire [7:0] index_addr;
assign index_addr = PHT_we ? PHT_wr_index : PHT_rd_index;

simple_port_lutram #(
    .SIZE(PHT_NUMS),
    .DATA_WIDTH(DATA_WIDTH)
) PHT_ram_data(
    .clka(clk),
    .rsta(reset),

    //写端口
    .ena(1'b1),
    .wea(PHT_we),
    .addra(index_addr),
    .dina(PHT_wr_data),
    .douta(PHT_rd_data)
);

endmodule